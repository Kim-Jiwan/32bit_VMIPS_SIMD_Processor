module vmips_top #(
    parameter instr_width  =  32
) (
    input   clk,
    input   rst,
    input   [instr_width-1:0]   instr
);
    
    wire 

endmodule